library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.chacc_pkg.all;

entity reference_processor is
    generic (dInitFile : string := "d_memory_lab4.mif";
             iInitFile : string := "i_memory_lab4.mif");
    port(
        clk                : in  std_logic;
        resetn             : in  std_logic;
        master_load_enable : in  std_logic;
        extIn              : in  std_logic_vector(7 downto 0);
        inValid            : in  std_logic;
        outReady           : in  std_logic;
        pc2seg             : out std_logic_vector(7 downto 0);
        imDataOut2seg      : out std_logic_vector(11 downto 0);
        dmDataOut2seg      : out std_logic_vector(7 downto 0);
        aluOut2seg         : out STD_LOGIC_VECTOR(7 downto 0);
        acc2seg            : out std_logic_vector(7 downto 0);
        busOut2seg         : out std_logic_vector(7 downto 0);
        extOut             : out std_logic_vector(7 downto 0);
        inReady            : out std_logic;
        outValid           : out std_logic
    );
end reference_processor;
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "ModelSim" , encrypt_agent_info = "2020.1"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lk4qQz2oJOBhDpUNrPoGwfMClfawqlxd9oXe2FUWHKSIQqQvSKuuENLEseNH8TWk
g0NP8ElUlHIXrDP76mHsRmavtir2fZokdSpNbjeE+9z+kOK/ZGbhOVBVwcJXvfzZ
JG6GFbasYNfJnRh7KluiLm2QtVhahEagAua/q9hJKIPQTBvJRpVUetreVJYUSIhI
10edhYWiU0HQE4cgwxLgCdHy7Qf2V0qVNfqDvcz0MKh+shJDL213ioLmZbDhKRNr
BdAsXKcb17q0eSQkTW/s0bhv3s5YdSwpSC8B/YIrbOyz13cNwagdjTtFmESo2moj
KM1gF73qH5i5MpMEJP+H+Q==
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 17664 )
`protect data_block
UUpEhjZxNiL2GMaewVIhmlljVwZWIrJyz2lEXqvEzjWB0QpJKb+9d7xDCh+ioQGw
rvg82dzcqkaRTNLFiFqpWhytuOezliHgCitD1n9rJR1amljMZsJAkO/dhudPsYO5
V4CWaK8mnH7xKXYdc0zM/ohxtLg1tQgCUzWRyxVGry0ogTuDDT4Pliym7azKvlPD
9ZGSpqaClJJmcgXZUqMR4FO/rUI+IgpPcp/1czi40jRtUQcLbgaazSKEzLTLDKo2
Cb2J/nW84S3l3LrUqoPTLsteRkUxShs/aamk61yx+H+ULy8+mmvb9Ehi46GzOh/l
1zuMA2XyIZC4c9yj1lLJleHMOSEowvviejOHda0r24FJCWOgWjnxImVqDEk3f+Ml
flZF1RUbcpqM35VD1pEvBxgfIDQVlFeNv3SJPyWBucJDfam+wjYPAe8BFLkkNXGl
E60Do7SQlxctbfPic1U359T3POTu74b2YznYUzvmpZ4yJPUbRuFvTa39gkMiLny1
MljnuEw0hnZS4ezdFKPWSA1bLQuikVuYLI9TOMpZh2UIwk8nnJMN122isPYF4w71
NPX9nTD6/shoYVyAz6uSet95eQ9NCjITV9FNiLg9B1lRNRP9jyVcPUAQJVsMNlQN
fdmL85KGjq7AeorVrJF1D4FbcKsrBRzDxOnFGsajUJvPRTyr+zo6T8tDiP3rZHRa
V/c6ReB5+SCqmARmq73BQymU7D5/D9r+4+Pq9Zluh16PGGDenRsQr/S0/pABX7rw
tsav/IjetplnZPg6tlpnKV4iYh+Pw5YDL54YZb6ZBoaZWPvYNdB5hs7mbEQtcX8E
7y+YcsZ6zFNDYj+NvtXlWM3+WDqS42tZXed7BVTwZhgBQ9RbPlCgMUFCUfEOSVw+
qwcIKtiENdtkhkMQZDJibt6rOWUIcZYyavlnJ38kp6V+oYjDbKdb46XiUyWWhFD2
sv9qkIbK2wRqXc429fsJJZk1WMdfRCwPvJ1dc5UKpHZyD707wxmMcbwF5pZo0lbA
fZ1KC22mj/XwqxO5PF7II26e1fBJm6BNyHg99sVCPqudF2DDnf/sE99HJOPU2Eel
7HIRdi2HH7FUwZV41kZvFpjK7QkRm5s3Dc3FBUAvb1PouSMh8Wm7tniGou8+IQOK
YHmGMWUUwvFBU3LJlfOKxgZf9wStBEtDTbC9zMGsh2uTls8xzoWy5p7tYN8z7+n1
cMSp91ItyvY9aLY+b4qNjE0O6A5dyRZYfvvxuSb56Fmu1EEmgqUUAwsNpyyitfVF
e4HNMcSkxX8JQyrFmg6PxF9xlOMd3clqjNICA+4pka31wR9yMyPcn1s+VIcljiVm
XfbZZSnFXL3yn4lH8mKb+I+Q6eVPXiZbTKACy3JuRzFW5DwO1lH4CXU/Qz4LcOIi
R9+AMWNVpuzPJ0uoy6GCH1YpzsKtww3ozjNEo3ifWjIYSTS1LJR+ITAj+2+GOqKb
toCe6UTeHddc6wiQMVcxbmEU5GGp4ugdvBxHjig2o8s/MH2U4L7MGf6TZBDWU+Hy
ipFZ0OXM6ZRqWwoWPH7dO78bDyXimce3fhBmw8rByte3QSLreab8lV/UFri8RZRu
MloUuxteFZqp93Pj3tbnv8PMmL6pNtUOuKISokzx8SJr4i5XSpxcVZ/Y9oPs09nu
wCJqrl92139SP7uiXWx3dni2CGqJMQrwiQDloKlgRMOhscRitltyecnyD2avg148
0Gu1ZJaP9jJKPtvvvwIbo2SPIsd3YMbt+tTWT6uKSny9kQBTDlKeSDcuZDkR3DI1
e6O7DYXgM8MeBkOdtaI63T19wVl9wTjRjIZJ0ZhS+aJWFkQA1e1ZshgI9CyIjV0o
EVrzAeAefavffHhu7p3S9mkIQ4lwIEO4I6WKXN5/dIpNtvhyn0WVrzt3HozOGP7X
y/EsWdT8J2qubf1oiRDF3AmInM8fI0Et/ZmFakyfdh7MA0I/gLuxCk8FvKR4mmBi
IPlB9lXX70qfIFgoHryXLq8saIl8QcI40bb0yO3Hhwff4pKZYnDIROtHe5FOEMvo
Hh0bF2UJjU5y10sLXM40UaJ/Vqy1t0WYTXOEG2s/7p2a83zhWOcRu1WruNi20pdy
NgsNOOM00UhauQgwHeavyHkUD84bC3q5I5qUZaKsd95fxkSfC7BkFNSUJIqh7y2f
1tcfajWxFIQ/8rj+uAobFXFvHbvnDaX8jzMH0c6n4e+5dUQ26Xg8w7stnGN2Bxhc
qOuQg2r9tzH5S8aYkDmGU5uLV4FjOXMO9y0RGI751HWae/pl4M8QufxjVwNXf3Ph
ZVxjmNwsj4f7KrqTqWAg8TwRhcI6tU0ECnlcwo9486ZzpfpYV+YuzrDR5O3Dm7Q9
rjd1VWEcHQaVHqpO8MLJL9tWUGih1arXF0i2Bb6FAxxptwaVhyFGYtTPrZC2nPmu
XThn5nxvLjEBE94uZgkiz+g3ZrvwYaS36+Z3U9/kjxartg7mxvUw/9laIQK0zrhD
Vnu8/PzPyQ1GhSwB8WGd8rWJFeaSzZC2OrtVkS0r6y9u5Sn/XYhpeHJPYur0Tvwq
He7pZh796sCmjSZAAgyuNOizgcq8aJdOV/PRBwxWWvJ3G9z8E0ShmdmOHzZDwc4t
7QpwmVDbQiU9whtvpM0a+DUyyiWnbMdwG5T0ch5QG83tOvEoLy4eIyUvJE+euM3m
xB2D1lvN1KEBjN8sm4FTW8Z4sUQDpxFjCUTlWds5R/uYtlUClOrsZUNG2tPLsqJt
rVxmI28+2flo5pw65Y4ee7O1XbX7LJ8XZ1h6CmFPBxx0aEq5ShccsrgMJ2nfGEvL
0q7fBsK2+HTq148psjl/+LJ9Py42ZgJCe9kwkV3QSbmIcasPGYtgSe0fEz7HuvEI
Nwroq5YICQQbLmDve9hWhz3pwD3sG1a+p2cLTM1m0dQzh140FUrZ7vE9VurmD2Yl
xeDc0jNbuN9JcKdk+5CJ9yomHeNXZNWjMpXhFxPSK2N4XiZWjK0qFB/bw8i5qFoM
MWN7waMcItz2omdy4sQhbrWdbH5NZFuYxyrAt8uq70oGltwmksuWs64yVy7sfMKZ
8uW+oINfXLJzq896U4Ug5+YKyX0vgOVkMiAxLrCODni3iN1TDWYkqTpBkDsM85iT
/6vukU5T+71b5AXIZWFfcOv+7wajL9t6ATedviiO52XWfbMPT7LQtW/pIdB6aJ4D
q68YxowItx+qxqYW4NYGmuhi6vLlbz2fIFijBzCkSJ4gPXMmBXJIlRuF455z81uw
rNkj2hye7Xp03MGhKZboYGvpjrJtV+MsIXHPO8uSH1oc0LrI3N4fgR3ATyzvfo2S
kseXrgZHs8p0WhXltV/4u8HGb6Y9H2FQQRPBB1bhZfGdYlYpNjbWqFoV6gRb1+1g
LzNYGNg4SNV1N46oUwl5I1aU8Pgq6MjmQ9I4bIfgLroRCBBM/QetZdU1cvZjvDKw
dJgZbmnh3ggluOuBk30CdHvdVXG2rrQx6fPMjtGoWugMX+CYiRYq7tdaYRmPpgnX
TzeGNCfeMxDjnAPInLZjEl0GTi2JnCV8MCa7KtN/xyDMsLm4IOsw01yE9MNV9pzE
oSwdKTAAMMMgWi5tfcsWrjUDIEXC3KzHfxDqEmfNMDG4fO3OscogLk5aB0TGQoQk
yQgOkig46gLJRT59ebMYKbD6JsFwZexVpJfRehIczpdlWask9Ed7bjG26LB0YICD
sDZQnus6cFrLl3IepyAzvi588RuY37azfJNFwUEE2UMHqVPAzzFBn4sozHs6D5/d
lGrA+uOXYw62AJ/+VdiOE3d5smjFyRhVSZSEHLDG7x2MRbM6pRvtZ08h281GzgjY
QMhGqyejhgWO7sSuWq5qe9ueirkm3UUVGNMc42d3bUDQYeqR6DAyvcx1a65QEpZE
Tezf9HiUs4BzJPmPCOHfMEy/sYdML426TcpZ4F+9uNmEDjjDcw2Rw/RzgRy0p72/
cX5nfVZNIm60dvKGqnYxmi7itgITPWVj8H80MKYVXCp4b8x5Y1gcxqL2k3A3BaH3
lXwJnaEDUNvjHCH6y5pDDqYSCyVGRiVXbrQ4cU/KzEbtYaahN5nUixZY/XsnNX+d
lV8I2SbJF8pOa8o8354w7m+vz5KUJ9mar57ce4e7IAUfKoCU1SGv+Doe2QAgXF76
O1PeuUamXEkuvSHdGW/pM9+a+FmpMHCGl3rvWHSz2HBRi0g3S6zM1PI4GaKWGlqx
CdyKr1AL6ZtA0JbrATwnA2JIaynx15clqZ6oX2jGYXUTWQ0plXydMkHwKKyUJKiM
Sx0l0A71uRUuVQAAxwgBlRLwgAbejL/gSZTS12DwVf2V0Pw0f+iSJH5Ot9RXFMUQ
6YBUPUgjE6sgDLzoBnqyO0UBc8tzSQ8cJb509Yd0pYcXDaEjVzcKsUAidabAj90H
RsB+VquxP9ZQ/bAPZ6FtVS52ZROBMzo5t6miexiyniuuN3OCxDEvmW/vElUkJI/P
XT/lcxWC3eO2HPcynLQfzIQhwMJg14qcPEZ8xew4qjnlZSOUgeE0b4RPD0OhtyY0
vJdsw8YnosVrAoe6f58C7X0rTJq4eNkNuzlJtRVzhpyBH1b7UdwijcwoVVx1VWV+
rnXJvX+hSAb4xcnTJ23U+FerPjjQCzJh7Z852ArsxUyxsSzvGLXxSiWSDBIsIJ6y
7dfoE4lGFjOngqEoZK9OkuCctOTwOa/G6tpYUOhgUu3ucT8d5pYPig6wIIKW6vwY
P19fk77KvzBtGI1MnFHYlxbKJlJ4PxG1S6L5lHhyqVT5MYHCe3Ew8JG4dbj3kWU5
gdQ69KEzJXdUNZnYt/FrzQfncahFYSbMFGVmZ+ZhKc0OoSRcKl/bYcB4xR+axaEL
2RYGtN3pvBkIEsYRY7TVzHXMldjibD+kxPNZ6qWcjb9dEhrRXtTAY8HnM2P19yQv
E2Act9Aq17mMBZhuuFSPt+h0EHPulQOX3xIradw7QC1CEVErz7xBkusxn+jTcKRO
aPqUwISGfj7YZFInjr2G0ejsa2A9FzacXU0a7TCqdcRd+lHfBeMI8jISuUH3uh1p
FQlG2G35XnvfBmp7wV4RZDZipDLUEbsvIkg3SR4QLjhjmZwGKpBk6x8XDQV8L0Xs
QYgrqVo14G9DO0rNFr8KLewu65SAg+p48S9/JNsBqSxq1RhBE/LV22JMbKCFRpBr
IF6WyyBdN94595ebNkOiREBhVp/CP4Fb27GyZKU2As4TzmuoUj2BhUXDsXuuigFG
Wx/XTd3lsUQZobP6T+KJOCmmYjE0TKOBlkBcBN1Ax5JOQGyKFsh+U57l+Dy1wDw3
rLZZOIRHqskQrls6bS2Sj5Ntkn/7CnMBTWqHA7UGFBCSTl+gZ/m8s2JKIVF/VIbh
jhgHANK9eg0QXVM6lj2sSLDgQNt+7syx6CNduuRjh4L121Zat5qVOBXk+HYvZQAl
m3i6GWW0tGn8QqBMwRo5ynnmcOMDfa164c3jTnMbWq094Tz9IZtFepJVkdU8EmA4
nC6cnxO2i2kc3GQgYNQWr7UIwLaxZs4u9pB77eXHj/+WF864HCyLRg0w+vr3kfNs
h1rr+SfPzPlmq7xvAXv9+cqN+toM/uy3w+r4LJJzzsLOB7ArI66Dwl/KJLVH9ska
ORkYM5LqoCDFyY7kTduyGsM8HFp4P5BTNl8QihEaZN4qKfCk6AUF3O+sdNCmzLnP
CsfsckXsbcxdnJoH/J6zaD36t5k+2+P774KORhM3/z9AzmywcjZ/ahRyWYS7KGAo
Bf6EJHJOS7xe3zr6Yr77F58Y06gc9vfkmCT5qNjXKHO2ycz1AIuz1ColL9TQQ7XD
rRLyHGzyV6RDuG2PhJDCQXufUVQ6gtaWZxyicZVYdukXSzu7BhOmiX+/XqXg9lGH
GHTDvm6OvBFsktiRBUPUZZS1hrNEsj310kCbX8ydH9VstrLxM7RUhav/jU79GHbc
9RH2btks1D9xB8bv4hTpB3ZLn3DyS6K/w1UE6vCGSuhDvZaa1nMqMBBdRuGpxfG6
SYR+cmHgoyakJI+S6kpdWY9WScRU67ntlRnbaL53LNE6hv24HNDFCscB/a9e9BGr
YEfq9h69ZrTsP4lcTESw1E3PuwTjaZjZnf/BkobxXZOpYU6DEtqGxNzWTUJiXD2Q
xVODk58F7hx1ShFVOaGaFEiQPkIdC3+Kmur7SBHb1HJuXNsFMVfpxdkllui0kXUS
arevCV9k4uqppvncggd+Fp2xJ0xfgea7ktgMAnw1TkU9NwMa//NOGLGXt+LDM7Xu
M765JOxFoylTZ3fL4EPAG+wTO1bb+KukfAGiQj/iQSZplShSVIQJvR/3gvUD3T/S
V5zvbTrgYPQgx2pWfIT8GDxXBpbq03o2jwIcH3Wt+DCh6smJSdW8Pp6kBeQ2WWXZ
be9mrO2KuIpSZJgUNgz6imKtvu+RtThEW1JQvtMtuiu7ZT2SibWxIBBUqyk0I26a
YAMU2m843YTerYDNB6hELtDaO2nfnv1+St73GykRm56QcsCSog/pRapfnF2PDVz/
Lfh3PXwvaLLnJCc537Xg1piDbNc5CW/WeH7wBIrC2Gmmc75A7zYZgvfrzDPCmyY1
xIxoTb5037paICpj8N4uw/q8KO2QzTlWgic7RxAxH84boo+7PlTrq8pMWUUi3QBo
h1VV0Gt/MQC5F8uxmXv78bayp29TANFr0y++Jq3Z3XqqLcQnkqLRZGHi45n5tO8C
kZUhvbLUopDlNJNJeYVHrJ9bf+vpsI51pts97O5Kd80gIZsxhQ0YWxuuVYJp4Ta4
jG9yEcRvRcQBB4JQIMINEkes704wmMq5mEXZID5PXrSioHAIwDgHmLWwYH0uWD5O
1/zLqtMtdZkKdbh1a3Z0fkmRSMcRGPUD3KRh6/Bk/xBdYkIaxvZg0c1NUZ+aN7B9
VCyKfRYqxzDXn610CgCm8Y5ira0vNgBhikVVIuAR5oW21ndH9zntZ6kF2DHoiavg
8RI3oiLKMrTyYFKqC2ejui4Z1eVGwKsvDxwgquQ29kAwmkG5ZJDlhw8mxHpi2nI6
FxlmwfSzmvRSwJFeZaahN2Kcy7v+qdv44vZ6nJn09KZ91w4ET0pt072oQbZUjL9Y
7LYI3te6GiZOFIRqCEtdBEu0v5OxG3pbM1qTFWZsqYGT1pkzIK3Sywap2zTq3Dhz
G5tkjWClFXWFE70qlQxEN5AbCEnRnVRq066tdDIY4A0jIbdgIlhV596DMEZ0PlTN
ruMA5pnYJESUv8sTBf3uT0mUhYZBpjA11+nNIZ99a102D4MX4xMXtWRIM2mdhqtz
WbAGZb7enGNCmhFB7VsN/UxJLmo/kfIPyclm9yxOO/BPqgKh+PyR19PMAQXAno9S
MNakv8Ik+UHMSerkkYFDH1DpdRHQvzeXyy0IjhHTpi/ztbejK2EeYmwyDKVb9PbG
Yxa+NKR1B39IFL48FQiIryUDRdviayNasV4R6iY1tBRqhdPSEFnNC4GZlgvjzgpT
Owt+ugcjM5WoDo3x38Zw6Y1E21TcBsv/i1mQ/x0IQ8kgJ0kdeksN61AultdYKQ99
0zX12cNMP5c+KuYPrJrlGsKcVBPe9rGUCey0egsnXdai0mMMoDP7pThU9ryEzihX
isDqPh9XJ6ce1LTMIWRQY8WdtXOZh0xhzTbOuMzdHqpnwuLJEKkoGL7w4HNKPrd0
KcmmPw8oyGhfU91jXVUoQIy3bNNmDCZSoHhclgoLFjcWbGlLeetaSSvfzgB/UiFm
dhkugECy79mbRCn5fUFC1rRjFEFxdOyPkvoGM4rW5Rwn8xJ/l5TK5zd8gAHpaf4L
tB5KcQ4UaITmAeQwGU1g64dBMTBQcNejrHQ5BrVNuPmvtEO0JZzeXd8KHTX7ImpO
XSVnsZmA/nHk5kMxjiilEZhncLPgSewmemTX1Tp2va56IHzhUHWo1ItEiN+cWLeF
qwi6h4LDrrOPrcSlAdF+xFgYrnuD9KiOZfgZg1lvffadatSxK3proBAMpUQzPKz2
bAmx27iUtqdEiYv/eSdifx5rxH4JWawiwZvCcNdfsHbn4l+SZWvO98BC7StXnzFr
RYt3SCl4uMJ51luehizEjSgtpNWFNXKqHhfWeHHT+A9egtIYvo5KLvgypZd1kpsE
wRl4KgK4tP6IOyGyV/iw8dpQoexIOH+4DiRUQKSWQJGLr2EYodUJ7UOpMzBgUjYp
jP8INdo5NSBbA846P7D3gAkmMfsX8GrMirvTjTW7Va8iG82JrfdgrKnowO7m/Gs+
CuFJpVF4mWlwGCEaEVfdX6NXABpY6pKRYZoA4XAtRB0CFvi1RoDvo2zmPNSabKjD
oLUUJUmv9/KEw60j3buUhW+C0wuq3X/Cr5PrID8TMbV4+g5AZwy5Cs1aRZRZUziW
q/klwJwqQ6PbI8AhBJ9lw2FRjpJQFnjIcog0X8DTzP0g7y2EEinOvbzACGIviKZf
VQ/xvarEWbcdVAfNg3rOxwYh/FmljGG2jTJfUZRjSTbsYG3dKYMeZeTgL+kPZkDM
Y+c5t5pGHb29V836stRzeHFLawkE4xJ+RjbyNeLIdnErTqgPY9+MS7Kc5u4PfBG2
0ECQt8y4JOdG0pMmghjO8DxVO99tG0IxodvPgASdJmIhHOE2vKmD4V464umZC1T6
XFlNFiQKOvu2+rLugiI+WTCWX5sBcHbXbv3UIhjAdO0Mx9Wh662JA1+jieSZJmA1
TTG5II9MeRAZprYEmKr5Z5PO3ABuK6kzfADoXQ588k7H12ApsXTv60afkAmx4Acs
N2D7mFvzRBLD/tO15homUNWMeSxXfxP6PwPeT5Pq4xQFy3lHUkIB4uHBMg46L3iP
XutGjNFz2M297uo2WRIr98e99RI8uILxlNxyP335uooawPy6eYNFmv+uZe3E3GiG
9hixDyAsio+cv8YNwbrpvxHFy5M2OdIYWbNijSXnbPvbycRxBKcuqJzBdB+J3ZT0
EJ6DbZAva3dNXHlBCKMwvSquM7JkIbwHY9ToHlksZjWKg8DXXP4AN86lg8tAXB9T
X5o6ROpTN365X+DeEyJDagF9DYlDkhrWaqVnw0BPUfUcFxg0OFteBV3OqCGv0MEN
dIhLvNawLKc+snGbNN8GX/P8Q5STChUjwzgBYDm0qVkClZfQeO+1ipaoGTIpzIqZ
As6mHRtyrSCq2OLiYWwU1SY/es3Yp8hrFA0HCb3n938uo7ui4RD35LTfYptKYx1G
IMkNPfA+zFaulVjstNlsDICGJEmPnu/E3uBHMD5/Qpje0EhK58UiGn+oYuCSex43
Y+VHIgqBiIzB5uCk6mnoq6mE4R610PWCJdkNySuViUh5Uhli8wzx84CtLYE05NhN
CqCgH9e5CNb+55FcZTN8VQ5Olr5ZStwSoN6C3PR49F9mEyLLW6O8ovAuKX+bFoNm
f9PMUyrrqkw1xNvwPtbhjCaFcz3qqAemcmobgpDHDqz2GfnioneJVt9TQJKqHdw3
CXcBOtVUOsQNfhoJomOhZF423OWMbKkc1OZhSERzJ7VUhY+kvUszkhD4Gvvjiq+J
GnoNn1gJ/wP6eYlYeVSwNUH0mH+SZ8ZSBhs9SaXfH4pJ038FXek+TyqSm+rS/SqM
ZfzfeQJgWbsngvDPrU/fl1F+LNnu3a1GK5qcen56aie/kcMZURv0uOQrQC2daVKJ
7ZCbC5w0mw5u4Ws40M6p5rH+KktWzlTw4VvUSeMTWPsUQJCl44aR3ouEZWNE1Vyy
jM8B31bldnMQwJUemYKsJ3Jklx/Ssl3jcIyKRRxnyuE3DUf2Gv5RC21LJZFxgR71
u5VqSvnyG+ACexErjpAsomk5cT0Fz3oFtp7pBg3iJBG9+VOYn87V/YouU4/WInjf
HrbcaalTTCIxTkxWk0XDhMAEQtemltu14yTHlg7dSebxR8ALb39mhdEgyZaKXhEu
TdCMzxxJ9V8DyLwWL9IP9peeVBl5Nf2ZWUGSXqJUInW6V5RhiZ1ncf9FcSH/e36f
IpyT3nnjwHiKwWquyLlX+RD5yMGG+UZXenpv6Fer3pAPo/QNzKWjhZtuK6h3od2B
GgJxVS8UmJpsWGICv0tj+dFYp+QIktZqjwUgyFKdyIyYY3TAUAb1UGRGtRsh/KJ5
sLamPSLIy22aQlmDQ9wDXv6QSpKXJU4k2Pn8qg2yoFfpxczk29siv6B5oXhVQWas
uZvofPu1CmzSCtMDRIO4DgGraJhOKzzapSZHlRHCeuTmf/khqvXDMb3+o3SkVk6y
n0wcW/UPVywDITQZWvTpqLJOKiYDWm99ydl31dgc3IKKDBxLxCTHvrq4nduQ5KG5
yL0TuIzeUZ7tYMyFucY2RN+vqyCDxJv/l7R8nP1dTR0pohCRgxIGYNBrt4JmBusQ
5v25T/VVrhxlqlNGUQ4YtkYObAWrG5SiKi/Q8PZw2D8yURJAi18ocIWKiwMVaaju
LgJte/O5+xlkHTiQ5dOkC/gtKuo47LE/LKms6SzDkx3q6S8QbNNCfC5fY1nao327
iQjJJs7530qUXYBlkQJxnJoiI7RCUuwiFeyC81nV3O+/+vcx0lYwvoSHUynVXuO8
KxA8dqHr81KMhPlmMi5WsZzThfDtflRbs93dykWLk/welwFy0POEpgfelzO4TgLO
7DrqiGDkA5WMt06lBaKhERMtdXvnCVJIDV4mQMXtjXsAwNh4Y7zIDoNXNj1f7vth
t5qLgzmYN9v6Ct84NbQWsXV6uO87wvuur2iHEpFBf0XidBjgV0NHNovtdgLluk6B
/6fTqGYJzKIv08dYevZ5La6ebCxH1dIWm/PRA8SEKp7cyxBuSFjuSCu2CbLc64Pe
M0valQ7tiRxUDB1wk/5yiMlOwC90gbhzObKc5brLm6qwkqmjRxMBVH7dh/B3Q5M9
E816u1d6fvGhslOLjPEKHIdAFMnNxyRSr68BmShahkX7f2y5bJ2CoSWDNEgEmW/C
hp9RV1Ih1/c3Q8Y2/SuHpHA7XeJrTCYRgwi27ktGP1Qegott/jOaLzWSJbXT3os0
UzgU9e5ix5irOi/3YMj6obsrjW8Xb5aK2mRGBf8XRgPaSDwTqElo3SkRQ9nHotOw
x52k097ZJ5G2RsjDSfEl6ijwfVzZuQzPHO1IVoeifge1Mrf9GGvNOdet93J+iIjQ
fGdcBm1mvEjE65TuJ8cKuXnl109r2meM3ORIPz9f7BfVKz42aaTn4Pc4KH0jhYDK
5s+tl0PxxWS+oaQmRwW0s1oPpFTjPIfrdWeQUoTiJi70Yquwwi3DzjHsNaRo2PGn
KYHAxZiF6ITrVqLW0jlcR16K46u0ABFKQaw7lWkyb8BVFe2OLJgQrQ7jLrbSPd9s
/b92PFzzB/8/UDLL/GM/4RUCgaZlNbT6jXZtMFxMiNatGNoqU9smamcacsWpPSW7
ColCL+FvI2Llk6HgEbo2mg+6ozOwcuFBT+l+nkTV79l8wRajAiW3TXrbDqZNtLk3
XP3LZCTdb+2d+4+tUpsear7L/82bv73ssGrLKxZooA1aP94sXc/Eu5c1mmcKYsBd
+gBzSHPWiruvkCf/ji5isqt2hgKHYcuIFxzauLTw1UmwzrfrqCdT+ZsAke/v9avQ
yWo39DrwamE9mFifij/JCs8atUcWNVkmyexX+G0ytKp6ZQkBLyo8Tw/0pMrF5AqG
EJpgulNVuUQlZa2vA7rLgwlgRAQwTs9HC5gDAiZqF7Ot9Nm4a/LVAtJmjym6Krij
yuyJWW4Sb8XvrznIllx1tPsMaMcc0L5EScknKKJVHC3sEmcthol2GvBys6vEKYqT
1sKcVvaJEgTFnoUSKxcy6NUbJjOJmEdu4JhYTAMYAdf8XMrGWpyEvpd/bevEJDpQ
aa3leikwOjBbIUuEYwfM+DyYXJIbyiX7bvd9Fm1ixmr8if1NM3B0VgS6glalkQiq
vIIi0Krq9srskCnNde9DYxO2UkRgLa1BBIlMRjuUiMeWyiguiy2B7u4zDIBGpNjN
/22EzQiFE/R0q1znq8XqkN9qQ5U37ObT2LhWoKZrJTEknRmsuXHJf+kDEmm8tY7h
QJ/ZoVnT79bY0a5vQjmerg+pHnn5TandrbBo/BJT5mT8H6j3Pz3JRwAPorVVfgrv
8dYdgvCwEV6Gy0tcFJERockaHGg5mPPsXpiqDYUItjBxM/POf9uFLKlxYWgdkEg0
zNMMD1KFJzxrmEISAC++sCjbhAQlpE3f9coKpuM/6OuBKmBMVuwRM65l5lkaPUFI
5iLwt4ldYiq748IRpZbn11sNOI52knSDegLGyugXoioTdHbVEWDffCwcqz2lusOY
L3ie7IhxenqouVJF0XBCDSypjpdxGdlVAyF04KIOjV/kvZTtJLYGR8ggucQA3SiV
G9PrHrSKP7Byn9GTX2BcXGNhYRLols+fQnXsIJIbPnkz+Q9YEDH/WQfL9uBr9JrC
SHzbLRycvLvVE1qvQ0O+OJ/TMgbrLmBNA095ixNc/YUYud/W2SrODfNI7j2hbJJm
mJbMmP9iV0h0Xmazg2eotuHxG8HzNMWrtJyqKLNqUzGJRWAd/JxqOomuqQYN+Je0
xfIckts3XUjQeKiA1EXPzwwiVyQrUYCCSfFKt57Bvh+aBDrIelbAVfwduPEs/iDv
zJ2wVlI2SHHZPxC3OXXDUcwoq5qhRGhc2wV/mp4sYj1sQw5o/1ieFRFfvspFMYnb
/ODqcDwppG4KdL1JxNJ5xWB8mNxbv6FPdfF8K5Rjee6qfw7AByZlw17+C8d0hEKT
F4qQ71MesUULNRRHR/06iHOuv2fbnDzyDPdZYWaNBxN+fxAcTC6uCb5N9HuTJ/Q2
zG3z9LsDO9vPqXcyPmYVVX1C1x9cEUeax2fKSVFuP6rAVWpu2URvT7HTd4Qk1mag
54T41b8cUZ1cxVMrjVKFgYyJqxN5pRiRH++5ExC2eJJeVF+lV6yk7Cx9/mkILmMD
JlvCOD/IMsB7Hle1nuoLwq4ulFYzSmSaZ8cS4oNxBVN5k/0lsxVDmFPnEgz/lzkN
qyjsjPW/w8fM4dcygwj80gKWAdUgp2a/bcooTS9SFGDA9rhZJ4lsi7TRZ4J9msDr
qQD0niV8E+wzTL0laIW9tXWcs8gbQq+J/Bvf/3pNPY1nRbpwFXa4g79ZfIgtgu/i
UdctYwrvoV3HPiYG/7a86QCB6jpPrv3WuxreEO4XurXR7FSW08AFpJnmkfP2/uPk
aj7KjGAe+rZ+vUczInmeVaUjrO+1xIppF4JncJI9Ef1yqWpKwoAF0N6hmrCTVR0M
s8IPYRqr2cDjuqMu6nSVjMfxQwg8gnLk1Rbh4AChkEaR52mI3cJeqFis+4euvv1l
C8LN+F7Z9pQquqnIYJ1JPqx79pyhh6rlc6pP1cf24Hvt6WeC/xZDzuvIE0VuvfOe
dZS42JqMs21a6n5C7U/f8u8SiYkW7qbOKgrL1GpUNxHDO9GpKzA6LSuBhRGSf2jn
DoewXWPQ9SqV14YlgerhgM2AwCgyi27TITgLJ/zVo6ru2BAQpPw0yN70PYe9vRDm
6JzAX6ZZnePVyJBfxR9GyG1t95FFg5HEiA4Y3cCt+J55/7jlJiUFFdsA6y9KqR3G
dLVIu4d+hmGtyyR1oqJNu8gP0HxiPx5kcEkVZdgMt03Q8HwVbc4GAWb2VmJoScyS
lG1AS5rbEB2zDKxeFrskBc+AEW7ojhk289iyG6kJWaCe/PcYkoCCtOCCdd+ziuAm
d+0xNdH2hzy5eAAUGGZKYDLiBIjxgrKUhCSvfwTLzbhOVFUVhIM2j9W0yxS52RCb
wJrU1gwxaMk6k30BFZQTpLw101ZNvX+jiHOVotHsE7qQZtt3vO68aQiZ0t6U+lyl
LfwziAgAIr62LC2xKa6Ov3OvyW3mu62+rcMF/CRXjBvRr2hciVa8r/T5ZYqY5aHH
0D3zptPQbrJf9+a16N6dVc9w7pHtUp2IvZ7xWGXDy3dJN06qBaoxs9W4P0Bjye9t
5WNRdrXVY37tu7+1MID/AfCciKlcwnuCyha6i06ZkKvIpdY+NIB6GJYzPidMMQ6X
vFioLYrtOn9Tf6zqaNMj7J4DqZa0zmo5Ey8MNkKBhWz56AQhrjndzNza/ctEQ/c3
15zmu+q4W03j5c6u/DrPseXYkDsJtQB+ZEoSGjez7oqZAmu+ECi5PHuueN56vMTA
FQ9QTbtxlV0c+0BVcWv62aGI+s+mJPy2778g7EMZhJEs+evCygPKLuBat2BOHqWQ
SzaIiy7yA5JGjK3kpVOHknCgfZSbi23l/JdI7BbmrFTkESqKtpxQLfjEAWt3KbvG
iAA2hAr1w2aDhbc9Pnx0k3KYEX2pU3AT7VDqTqluZtVwqyY3LdI0/U1hj4LL/KUG
7ByXe+T6M06ynRMOJU/SeR5qXcxJcyevj1oqNqqRhc/BoUE9Y+3o8OR1m28uc4YW
Igde/AIP2GWLLz47ky/265zlnnYts8XXGA5X/eS7VOZlPh+urbRFvkzk5TbULoJA
LYUWZo1s3XhdAQWQ+a2Oa9LC7s69R9z2WLIwFQSU4lcnyrnTUiGZiM4/l8dbDCqJ
dsxaWJ8G6EhHlaDRfWhIEKtrdMMnjYElX+lldSUXWGVjfCnnQyy6Yic46FJB4HBK
lfmcpMG/V4puHiSd4qjcA89+f4js8JDOVdGQ/+D3DsEBVN2uO1qagxs+uqtpkMUg
ku9Br6EO4iJWvIOiwoDq0AXnuXoM7jSo4FxRONb6eLtk04mdUKJBD+8ZEAFqW4VD
PgoobtW+cMpN5Z7LIj0j3IubRKqGPxAtWHsuQVrnDwou4rlAor/rFJXYDOTd6jV0
U+Ad+wWv/jts58eHSw10uZSYUtaHVcqwn3mTLUr5svocofbzQg9fyVkfpfgQ7S9y
FilyJk3ghRUEazYQe11UGYM4aLQQIEhMq7pntaBy6i5cF5TfOEsJ0daP3rdWEQZH
1b99AFD3/LZnr+HGloTEDvgit0+YySH2ROS4IW6IkI1iItXbqqt5bQOuxlae/w1B
USBmoxqxoJwCcAnaUukWiPSgUsDd4UW8rRWb4EoKYqJYbhjBtph0cObkawyC/Gzh
vSkWyWV6CNImX8q0pXnfyLuMUr/Uaoglp3Xigp8WsCCaoBuJGXgwFQIoDs3H6oM2
ZCq2Qe0yWdw7X4BM+qVz9rjCpxuKhliVImpYrnCqEXlXV1CmFZzrgu7U/qc/LPaV
hGUMesAMECflHvTELiodGt73/AgnZbZxg/MauwIrsW1EWJSwGrqi6nTFuBe267vH
ygVlA1AViluyyDCOVwcLO2Ofkon775MEjhmkbRaB+cw+ODFhcPrvjolbXmlNpbQH
/wQnNTXOvuqG564YDfdTQ2NvSy0Oxh4S0hBiiY1uoLbrK6taIrq2CVmV9yUesHxb
UbYPyPJhcbfkGi0dwD1PV1vCkAz/N6FPIq0/Q/OCwhs77dJsbja1ow8aKEWM5eF2
FWCILEruMl/g08MiDPTPG9rXRPEeBeepMMm25U67/TMGRgWCHyNotXhOQ/2cA75b
VB7rIP53OeB80ds2QRbQ0O8bAPYeLylaTOS5fur4nBh7fX1HTpS+Rpiwv9XbZMli
5tRCnO0klq4jbfRQ79t3oMqXxBORLQ0o7TR1iBOJz35qNHqcasST4iN7c8DUE9yu
NJJPv3Aj4sy1lazCuECMq2Y19bUd4WMJJ7eune/+05Pc1JCjdfJxez0e1MbOI5qO
Ox4KMx41DCRa/mN1XpovmgtwR91EtPx9lw48DL+2lSwyHLa+R+wI1SqlnY1SLNEP
m+H8YyEdk+pGAXeLtJNS841pPnFXYY5ZT0fGQOrSWb2vvzjlANtDHtNYVnu+e/AQ
Mlu/yDocFHxT66iKs6pn/aAyEF1PUGxvWobk9v33x1FN31s2YvyVHGhm0KmREnkn
TggNK0vIkwbw/zspPZFBFhqn5hpOdiRKkVbYwX3Z+o63Oc3ShxY7HNZ3MY3Yj+BM
KID8XLtjr7ud36nmo3x0tghtVaTRQwFYh+C6PhW7S59ktzYvCL53u8YrkTc3jGVv
5Ns8e3sEYx3wibKOfZsI8zQA7i43HM094nw3tqBgatg38AV+00dM+qNBKLfP4HUP
WK5NBcZ7djMZ26UuvkRZCSRgNDIG1Y86ieGVEbXmAG1TQIlUOeB3pudCIddByU3C
B1tLPJcDF3tqJjq81ObUzJqrta2tP6A6FwCMgvhD2UZG6gU+BqacgFQrvKbPHH3X
ncm1EukN5roQACKfu+fHro7d8PdW37C3z2ngNEeEzuxOBZXWlIdBygV+3f85NNxa
MW1mvZB4kIIhNfVwnOCm0nJXtg+f/sNxz7WjIenP83i0MD9CkXdaVK+AAiDoLvsA
YFfBXVNqgZBlrW3a1HvwYZJdJwvNmiEwqSkAJryrxLzDYzwC9qTCuhP3nTkKLvcQ
aVC754F6ylZ+2W5J9/FZgS/za0nNi5a7J8oZ5sP/z8lW4+ehJ5YDubXbGNTpY27W
+qVOYg3YvTHbjHd6yHv919uuo65r3rp7R3ZlpQ8EhodIcb0CmmJGCdsixXyzNEza
5rlQtwVrAdzXTktho1DWAVmm0uVVZQT/ogafarYuam4zy2InPT4g1HK/wsb8fpv+
y5OnUORn8VRTuf7HxZfRUmXP7ZNkd4G3j2fQiPvILWb+aPcKN1JcqUtwGGZAaYyw
ERY8fbdJKhvueAF13vciWQSkv+71kh3YdaaUBhgQm/nDRE4qc1yZoURoXWiXfr9V
Rp6O6WJRmrHOIP9GJYgQZ2X5VPIVCpmUekFxAzrqbLLn1G0Cg3Zot3uHyGQxN1K5
x7bHiiuqELQRKRt/wH02AUP+qf16+wuRqysW8tgZbbpDVTkQmSxVgzwYyCqfBF7i
12T+rJIgqHAWhk4PM/TGRdAfZEbjbEoQOay6wXbDpfPhcCefHyIj8O+mK7e/Ar4B
6AydiNoiyjur2OMC3QThV8AzwFoYbQYAG4sNpFLDppVTw9Eh1uPaVUOmp+9tQLRe
rXCw5TQYunrnu5Ihx8caQ1yM12H8KXep8QoKfu47d+OgnrXcampybW59O1nXVYY0
Vh5THdLkEJor9mmx9fKgBmpepRuxwzMsuSUK18wC8j0cXZ3T3KlFELauP4ha4JTT
mKIpLxVqHQRlObq0jXEl9jMnEKlmdyZc/VMwPg+AE0zpSkUQbVYu2qApyIdZg5TO
mO88O5feRz6z1jYzoyPU3igOo/Wk2RIWY69IliJrlkLrepGkl0ka9G3IVpAhu0T8
vaDvIAEI/0X42ewYF6vP1OboGxvjp4NeeJBz2u+eei3ZchqBQsryNt+dMUkuIk3b
/XU+vkLEDljiiJrCBJC70N64yBXKjZIEskY9AclAFX5McpRJopHGMyq0jv1GG4Cs
Nqdx1udCFRCzYZFALTVIwoH3Nlk9SKht81HzrsZf/Od84hyfAjGk1cRnh7ZWMyYI
ZiPYerreLpJqqd8HcNul+Y36ApbKBe2Dey6AEDFDkXFYTpXhRvzOTsVFd/vMSj8+
lm+V83PLQV3nkJD/WfqC7IkctKYwoOJLlx2HxQpfDEL0AX0HicdkAbaQ8E2uGtkr
C3vRc80u4kjb+1kvG7fP1JFDkG/B413hQlAhW3Dib1oUcWc0fwEgMPidfk+R+Qc4
Erdri60KIlfPymn34eH66bt5v8lpVUBTZ5Rqo2RxVrFVLoXnkvAjAEQn4qyoycDR
YBoxoD2NRBy46OFnGTKI2tB714v8gXGkOCbJw74c0gCHWvPbpP1JQGDL5E94sMsX
9YaJprSQCO4mBCRiX2/q1IsJjgImAcgMhgj7H5nmxKzOUnesjNxwxxBSHEGUFSNo
EGEr76GWcW8vKTm6wx6inJBR1D388Btw4fP0HkWC2UiREe6eM2kMy7sBvmlhsPdS
4CtX5djbcmLvWIyXCyKQerQtNpzA77L8cAOfmX9EOl5689dvISsNirOgTcWpUuGG
VHFLm+7lx18PaUy8Gzb0mRInLBQXfdOUmWuatHorgrdPVeOpK9zsvSOuFuXkzuWF
gBcIc35nu8a6woG8V9H/NgIo8Ol18u48Oh0W4OKkaXacbvpxD3ONq2vBULbzZTh9
gxPNB2o6IyAZkcQeY1HLwXoWc0df8mnQZWgx7iaRXTrfpqGgBRaNqYtdGKO6+xSf
BGgV5pJaAfPq+dF9aLHJVIv+bwxFSR5IizYgbw16uXpmDKSxqNNj/cU69XuUZOZ4
hIwBHtzbVRkd5yjweYTb+YNRGP6Y9Nu4ec9FLa48QR2jWjaZ5p6VM3SVXrw1aDEj
062m0tBrDII/f+gtr3kE4VfeqTsmHS6+aTPGvWToBq2iHJY9f8Bp7hf+OK9d/mT0
Ifc2o8PcOJaqr4Lkz6WcWyT/ouQRlnyrrjKusE14vsH4jn1OLLPXxt+MyfwSKfKH
eXMd1RvXJ8t6FiCbb7NWthFxYbOLr2CudYqURLrNVwqOxHUgyTwqQGOv9og+JwJL
cIkcDJ9p854xmM4qBv/4uohCyQ6BSgiiztepFVR9pKqQ7jezMDqEivtn/mGBeKbe
ln9B/Icygax1bqVDLHRw7KrkGQZvtLUAdSLtLgUSSrFbw/RUvSoI55hAxApMU3LK
FnTeGD4M/3yj7q1/vZxUFPbUOMWdjLmtNWoY1RuvtLMcNBkoJy6XI/8g5CtifRfI
9Y/gu1IIKyicmxInpATxxPNXwB/yLd5xW+PPQZgZRMW5kNheEaQ5f8PKxU7+Z2AY
HSnpzGLCPbpkHfAl/sUrFKjbcEiHHpNkPetbM10umOR1dp3Vk/y4byumnykpJ2zS
c/jm7yleBMKnSmrpQAO18TVxC1pJL+uT+tk0qyBpih00WlhRQadf0leUX10ZAOlJ
gYtM2bzFzcl+rt4iESa/8DFaioArpfX0lRow7Awvfu2Ed5jGQrleVkZ4v87TdNfD
c4fYlGt0qwR4471KgZnKYDlCtACID4WvHQbkbDDJkXUvUpw3hmsB6g6xTuknXdap
/3AtY3ZgDWJ2iigaa8BRAy2TqTYT65/GCuqcI83OJJner2XZPfaJc/83lF+xFi7o
tdVMaLiG07UgOaMYrSVvnJCkJfvgrvOCLGPR0+MK+RU+KGcd+mV4dt0T74XUWcps
7x2peMETeSsQ6fFnexPxzC7Yj31Jo/jKDXRi0qSbG4yO3BbCF7TqC48dPDSreEfp
bKcboa9X6cOlpU0hFMyZnDKiuHVy44cAqCPHgp/bfZSRm15W4a5q7JxIW/tbTDsa
lxxzZ6p/jKaO3A3bONPdm4zebM1mE2v47CKJPwXPFQsvLxuNiPR4PFTt1DDbeTfY
FYENcFRkskd/67TpMs8AP3ZlwKQgKZ6eYxRY6ZNO6aeUfIBRVd1s6hTatmpxLaac
4Raxzm4JgQTOzvD7Fdbm4Ez2FyU1RYpvBiLwzZyZ2gn5ccHfdigQJUJpqu69qES8
2p7YHlBEAG2XIZwptZuoeGovkbFVmo3PgbWm9NSzpRi0BmJEo62/ucW7cj9wQSPx
ZFpQ54ubI6BOW1+mNuG40W0PTkP4FBzEyne7DorkhLr7Z0XDOT3xTWVVUdDALxsf
cd9xOL4hYeHuyCa9NYPcaYl+KTGNY/HmFAEco2UvOvEExyGqBFVOjKD8hQ5FCx+A
+eT+USlxwBub8ZP5rEFwRr+uc3S91Pp/rVtNTEPRWtBliHmVwV468rFubEbCF0PT
IAPd0awW2ONcBKL8NYfu4UHv+/C11scfUOk9tDIQvi/UrRkYYRg4p5fgqjzLw5Tj
zDNXvSA680Nz2jw1PB6hoMRZ+a5zRYuAUr+AVPD/tvTVqXLmjlRxYZZKk698nugk
L01Kid9+UHyHZluzzM3LdMG5uH7AkCQptUiSgCcOu24qCcH7Olq74kEbUWhgqo+w
F+LtkfXfNAeNo2XXzUHZ6gMJ4u2Mct5cu+BwCD2cumbCn3u1cmSsC2lbu8yMWMcw
D+JmvqSL9bfJ/qqy+TTFMH4/OOyWybBfOGpylpLtLedHqj6ipPTeRRsZlGxAThCj
7PWSEUYPX8Ycg3K+SUR463+bDGiwaYg+qeparq7azOBRgxN9JUz5vHU7u3wTaEJj
PcMFJ9vZ/4IStszujwRU1zzQ9q0ePSDVKiCSfgvesiwsj/kif0I4MQ7GkD06O4BM
iwxToWtFL8osuZ27LW3bHiNk58rpZjybEK6dxgQvigjs4zZZT+9g5nxEfuiF4EPl
Wcp1YwZpqU5Ox1QekL6m1nZCyOcTsP1MRp38Sdz/0KYCuLZm+XutqZwpMlDcXncq
Aro3SGovWIfA6ri73+oz14Pe5RPmITPVbqweSV66SNETJ7DMTkr0SMpgb6VkD+pB
jGDWPPgVcuNF/ujHzIocIiSzN0SNphM04B4LRcK9/9WGPYmNXFIhcGPalW5i+wl4
nogjSMlV3vBC5wIZ2goxOxSORFlpuwGY21M5T4a1XlE+TBWTdEmGlj0a1ae6EbeO
JHiT9QcngP0QJQerldsopMZ25zc40K0j30vA69vG57vuakFXoQUGxsgUUqgerKmp
wyVuQSAT7nNHOvrHpQVjqoeGk3MXioZ0lLKDxjVxPYV/wTsLXX95iupfk8Ic+ln6
RHTtuxvqhpvlXgOt1nLwINVr1+EzBMAQXh5SfIJ8xBlW8Nj+BDYnKPUr5nuEOvnV
dpnPCu/9lcyTyRVo9KQ7h8yrNQxR9kCTU3Sbc+VrFuiTpp0fDzFZ+oxpeNi6B42+
JvDAvtMJeybXaHugXYz/zjcjcCKb5l9VcqlAYHrDOgszfn/Z+B8khFB9080zx4h5
yMIJfdZ8WO8FbOi7boGZYGaUGRxMj11iBxs0SgubMLt5R6Z0aZdsa0rhV3+cAhmZ
jhjIpWvsfvpX3TIfo9g/ZPsgCzBjd8RKn55dugdjS7MuBtezCKweCmJQZglYo4cL
RLfNrMXx+GraQLKDWMyq6BtdEPZzzYpjItlBfIhWdGNIEsJHcPeP291JHa/fFdrg
BdcCOysqEZ3vxl6hoKzYznczltMdG2p22xrVNbvfNAjeFOV4qIvlZexZ6O9kyekm
RLqVZmszAiMwdyfQzz9k/M3Vg6L2HWGMJkOGax8HLc32JWCVc8I1/IMV7sHgO2gt
QBsMTj4xJIJJBpvdGizdKyFNMA6+GJd7r37/ZJ9lNgFTELQmPgGzxrp0NyvOanl/
UHMQKGyDsLHmyaJBfwmjeAB2Yi5meBautS7aU3/xYnY1gN7E2NxTTokXnrIF70gI
ba+GUhEtHkYA9qowivxXQ9tdW81YJdtfwatkbBz4ybeDt/ghFUuEVI4664gElQLM
7sCDceQsSPJ2QXneBItL3N9eNjruRwTkXGEfwx37XId09Y92YW8+UMvnQUDYch88
mMXHYV30mqicNX+utdw1R6DNin6FIxNRzNEFP/zhAIia2Kn/r/TpbZusRpin5iZS
bUuGltvv6sj+hOpufZLaJz4D6eOSsG5/fJHeaoVdfF4JnDX3RAte+9Z8IoEaD40C
/bueZiUeigC9XOS15fhrA3RBbycfPkhxRGO6qkmUbh0vhoiZnIPSBc3tmNfBph2f
9irWD39MEvk10vsFbkRZov8AtjnLfd80xlNmJoZuaT/JjilebYpmpH61ohn0v0Me
LE681L7n79wjIg4xfZUjf3R+/3izwgV97ovI4MmUBZWhnxe2fNTvGLD+s1Tny1B7
axHiq7MFioOKkqqp9mS0kREm49Xz16ZuQSEWn81nmx6xMTt84QKAiQJwzku6NJVV
+n0jZolcW1+yKaICMW06ndEZmRq8/z8jhov/P1lgi5Gw/bcxQI/Wkq4ezkMcGZ7r
KLycwmm9zlcaHuQdTy/Kn/VZCkjX+uX7xR4zcHzh/455W75j8AE/vgfkwCSyPCVV
XibP41eOp0iQlTW/iSHuZwsSjbL672ElfXvIDTd/CofrV1A5fe0OGS4QtmTpcMNm
0i0iHGbKH81J3dpf5JuJ8TJlWlAtg1NswQ7hGN/ZwtzaO7gISgfe0q3/bUvZIfVj
zOULhUNtCoGsaAXbfnAMWEIXm6B+yhS/3doIyjZmUOfG8GT+sceBhjY/TRtFW2p+
PLOco6Kr9waIv+UWhRgFaWnNqoMKhLrreENG9BJ/XkmS7OGtuJlk3tV+jAlnAfpB
xIgTqy+4UJRx92hTbo/F3jnoadPSVR2zrmcPIxsYSIAZGip736mOPYVkfdgNXZ3I
Nl8hBkyrrE0gXegj/6FNZ+AONF5l6ShqUMVLtbeMLY443Srpb1oF+wkCFnH0vUWX
mMZTrJkvqr41hywLDeByXmAcbUW4a9+NWE+tWb3e2xtGF3CgYUNk0b3eex8M7nPe
0fL6pnaZTiEntDL+B69lWSuAkzlTfHLHRNw/e+rJc9g3Lef7N79nnXdcmPqBE8BE
1VYQPRL0ztTKddwcBJGnPhKdGxMWjaJrK+O83H596KG7NN87ZcG3jZdb0jaIqULc
e5HeUfc1J9Aiuvjqf7CsH1EUDKnlQShVWwhCPDnwwlHr2iXDy6YLgquhEEQGb2OW
QMb0u3Clb2A35JUogVjGGFKAn/d2Ya+a6RmkbJCHEVSRmrImhqMafhzNqMN+CcAZ
9Jw0vBs6Cx7UdmbTLblnSo3eCWdfW+rfU68cr/zigzNJjC4V5g2jfSXf7nSjgj50
n3ux/EYUyOAsOFq3JImJUgnVdgRx2iJ0/IsJsRWp8DmQBnZWd9YyETCLMr20IwYI
6umzwG0Ay6Yt1POdiaOZvUG9ai+mhxiUMLsWE5W7LD1hGWdW4Dhua/74XLphm/MR
5ITx2JCUozR5ZKwo4Myyn4Uy0mZF4qbCEScZBVGWhlRmTNRm5CaZTu4jzzb9KqF5
QxTDqV9p/YVTn0LbWVFRrLJa9/ZUGCRbF20YjmveGAIW2BsCNobNZfxq2Im5pWpn
sqfUhyCGF5Cz3d8ezCNpKjs/tluDwy6SL2OqqcKYmL0DlcPgkLVi9T61m9PARvv1
RmdqDk+XGxoHnai9MVpRgTHNMFbx/hY/DZoJEnr+1TSdNUHH1n0UUssXmjbvVfcL
ngwEzmvaZi57bohNDbBUmGfrhXX0Yqe4Ma4J87xv8oSRt6gC3/XVEEhr4xXGDTTL
hC6HlR7Dm3glHOyviFJusyl5Ou7B0vvq2CZd/IJleeOMtvJ8Ta4cKfW99U4f4zTn
ZOhxzUbrtMqRQAMKBevtI0C16Wyx6h17zsild+sQ1bD2g3RDBRrjNd0umV937sRW
M0Vg4+1w1ObpUhsVdzpA1aP7xKFcY+zy72FwIYiKuDyH6n4fGYL7tj544y9BkWqt
4Akb7lnQKxElIUmncMRnELX7PJz8TJTMjWB++uI2de3EYDoJ73sSOTMbh31dX2cN
XOrX69jtRMJFeQ+fWcTitolg7N3YFWRGlQvWwVwz2qCbjkVDRIi/2afQ0FNFc5No
FFLNOvn1lA9nCWMIHR4sWDhdL4sdic/cmzoZIkbTB/llEglWvguxOO/xm7C35h8G
1Rxnn0yxnAosT9CiTrm/7XU7M+An7i6EgVZS4iXI4QpMfhtUtgT8HY2CuoqIeWj8
0+9E/ltXGcsP/fFiQd2qN/pQ+lBHBVu8dNAJneJCK79GdBPMdABm6VxjDxLDLJ0L
`protect end_protected
